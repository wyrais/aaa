module ALB (
    input  [7:0] R,      // ???????? R
    input  [7:0] S,      // ???????? S
    input        CI,     // ???? ????????
    input  [1:0] ALB_MI, // ??????? ???????????????
    output reg [7:0] F,  // ????????? ????????
    output       CO,     // ???????????
    output       ZO,     // ???????? ?????????
    output       NO,     // ????
    output       VO      // ????????????
);

    // ????????? ????? ??????????? ???? ?????????????
    wire [7:0] or_result   = R | S;
    wire [7:0] xor_result  = R ^ S;

    wire [8:0] add_result  = R + S + CI;            // 9 ??? ? ??? CO
    wire [8:0] sub_result  = S + (~R) + CI;         // S - R - 1 + CI (?????????? ?? ??????)

    // ??????
    assign CO = (ALB_MI == 2'b01) ? add_result[8] :
                (ALB_MI == 2'b10) ? sub_result[8] : 1'b0;

    assign ZO = (F == 8'b00000000);
    assign NO = F[7];
    assign VO = (ALB_MI == 2'b01) ?
                ((R[7] == S[7]) && (F[7] != R[7])) :
                (ALB_MI == 2'b10) ?
                ((S[7] != R[7]) && (F[7] != S[7])) :
                1'b0;

    // ????????????? ??? ?????? ??????????
    always @(*) begin
        case (ALB_MI)
            2'b00: F = or_result;
            2'b01: F = add_result[7:0];
            2'b10: F = sub_result[7:0];
            2'b11: F = xor_result;
            default: F = 8'b00000000;
        endcase
    end

endmodule

