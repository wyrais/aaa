`timescale 1ns / 1ps

module alb_tb;

    // ?????? ??????? ??? ALB
    wire [7:0] R;
    wire [7:0] S;
    wire       CI;
    wire [1:0] ALB_MI;

    // ??????? ??????? ? ALB
    wire [7:0] F;
    wire       CO, ZO, NO, VO;

    // ??????? ????????? ? ????????
    reg clk = 0;
    reg resetb = 0;

    // ????????? ?????????: 10 ?? ??????
    always #5 clk = ~clk;

    // ????????? ????????: ???????? ???????
    initial begin
        resetb = 0;
        #15 resetb = 1;
    end

    // ??????????? ?????? ALB
    ALB uut (
        .R(R),
        .S(S),
        .CI(CI),
        .ALB_MI(ALB_MI),
        .F(F),
        .CO(CO),
        .ZO(ZO),
        .NO(NO),
        .VO(VO)
    );

    // ??????????? ??????? (?????????? ????????)
    stimulus stim (
        .R(R),
        .S(S),
        .CI(CI),
        .ALB_MI(ALB_MI),
        .clk(clk),
        .resetb(resetb)
    );

    // ?????????? ???????????
    initial begin
        $display("Time\tALB_MI\tR\t\tS\t\tCI\tF\t\tCO ZO NO VO");
        $monitor("%0dns\t%b\t%b\t%b\t%b\t%b\t%b  %b  %b  %b",
                 $time, ALB_MI, R, S, CI, F, CO, ZO, NO, VO);
    end

endmodule

